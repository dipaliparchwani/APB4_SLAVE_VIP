module assertion;
endmodule

