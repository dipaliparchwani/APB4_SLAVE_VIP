class configure #(parameter int depth = 1024,width = 8);
	bit [width-1:0] memory [depth-1:0]; 

endclass
