package my_pkg;
   `include "../SV/apb_slave_config.sv"
   `include "../SV/apb_slave_transaction.sv"
   `include "testcase1.sv"
endpackage
