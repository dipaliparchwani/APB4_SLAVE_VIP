class coverage;
endclass

