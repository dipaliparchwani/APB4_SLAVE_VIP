package my_pkg;
   `define addr_width 32
   `define data_width 32
   `include "testcase1.sv"
endpackage
