package file_pkg;
  `include "apb_slave_config.sv"
  `include "apb_slave_transaction.sv"
  `include "apb_slave_generator.sv"
  `include "apb_slave_driver.sv"
  `include "apb_slave_monitor.sv"
  `include "slave_scoreboard.sv"
  `include "apb_slave_environment.sv"
endpackage



